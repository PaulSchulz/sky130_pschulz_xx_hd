magic
tech sky130A
timestamp 1598777367
<< metal1 >>
rect 15 75 30 90
rect 0 60 45 75
rect 15 0 30 60
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
