magic
tech sky130A
timestamp 1598787703
<< metal1 >>
rect 10 100 35 105
rect 5 95 40 100
rect 0 85 45 95
rect 0 75 15 85
rect 30 65 45 85
rect 25 60 45 65
rect 15 55 45 60
rect 10 50 40 55
rect 10 40 35 50
rect 5 0 40 25
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
