magic
tech sky130A
timestamp 1598785497
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
