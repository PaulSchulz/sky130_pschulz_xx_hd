magic
tech sky130A
timestamp 1598786254
<< metal1 >>
rect 0 75 30 105
rect 15 60 30 75
<< properties >>
string FIXED_BBOX 0 -30 45 105
<< end >>
