magic
tech sky130A
timestamp 1598838751
<< metal1 >>
rect 255 645 330 660
rect 120 600 165 615
rect 105 585 195 600
rect 240 585 345 645
rect 420 600 465 615
rect 390 585 480 600
rect 105 570 210 585
rect 225 570 360 585
rect 375 570 480 585
rect 105 555 480 570
rect 120 525 465 555
rect 135 510 450 525
rect 150 495 440 510
rect 135 480 255 495
rect 330 480 450 495
rect 75 465 240 480
rect 345 465 510 480
rect 45 390 225 465
rect 360 390 525 465
rect 75 375 240 390
rect 345 375 510 390
rect 135 360 255 375
rect 150 345 255 360
rect 330 360 450 375
rect 330 345 435 360
rect 135 330 240 345
rect 120 315 240 330
rect 345 330 450 345
rect 345 315 465 330
rect 120 300 225 315
rect 105 285 225 300
rect 360 305 465 315
rect 360 300 470 305
rect 360 285 480 300
rect 105 270 210 285
rect 375 270 480 285
rect 105 255 195 270
rect 390 255 480 270
rect 120 240 165 255
rect 420 240 465 255
rect 10 175 35 180
rect 70 175 95 180
rect 125 175 160 180
rect 180 175 215 180
rect 280 175 315 180
rect 340 175 365 180
rect 5 170 40 175
rect 65 170 100 175
rect 0 160 45 170
rect 0 125 15 160
rect 30 125 45 160
rect 0 115 45 125
rect 60 160 105 170
rect 60 125 75 160
rect 90 125 105 160
rect 60 115 105 125
rect 120 165 165 175
rect 120 150 135 165
rect 150 150 165 165
rect 120 140 165 150
rect 180 170 220 175
rect 275 170 315 175
rect 335 170 370 175
rect 180 160 225 170
rect 120 135 160 140
rect 120 120 135 135
rect 5 110 40 115
rect 60 110 100 115
rect 120 110 165 120
rect 10 105 35 110
rect 60 105 95 110
rect 125 105 165 110
rect 180 105 195 160
rect 210 105 225 160
rect 270 165 315 170
rect 270 150 290 165
rect 330 160 375 170
rect 270 145 305 150
rect 275 140 310 145
rect 280 135 315 140
rect 295 120 315 135
rect 270 115 315 120
rect 330 125 345 160
rect 360 125 375 160
rect 330 115 375 125
rect 390 125 405 180
rect 420 125 435 180
rect 390 115 435 125
rect 450 175 485 180
rect 520 175 545 180
rect 575 175 610 180
rect 450 170 490 175
rect 515 170 550 175
rect 450 160 495 170
rect 270 110 310 115
rect 335 110 370 115
rect 395 110 430 115
rect 270 105 305 110
rect 340 105 365 110
rect 400 105 425 110
rect 450 105 465 160
rect 480 150 495 160
rect 510 160 555 170
rect 510 125 525 160
rect 540 150 555 160
rect 570 165 615 175
rect 570 150 585 165
rect 600 150 615 165
rect 570 140 615 150
rect 570 135 610 140
rect 540 125 555 135
rect 510 115 555 125
rect 570 120 585 135
rect 515 110 550 115
rect 570 110 615 120
rect 520 105 545 110
rect 575 105 615 110
rect 60 75 75 105
rect 270 75 285 105
rect 60 70 95 75
rect 120 70 160 75
rect 180 70 215 75
rect 250 70 285 75
rect 60 65 100 70
rect 60 55 105 65
rect 120 60 165 70
rect 60 0 75 55
rect 90 0 105 55
rect 150 45 165 60
rect 120 30 165 45
rect 120 15 135 30
rect 150 15 165 30
rect 120 5 165 15
rect 125 0 165 5
rect 180 65 220 70
rect 245 65 285 70
rect 180 55 225 65
rect 180 0 195 55
rect 210 45 225 55
rect 240 55 285 65
rect 240 20 255 55
rect 270 20 285 55
rect 240 10 285 20
rect 300 20 315 75
rect 330 20 345 75
rect 360 20 375 75
rect 390 70 430 75
rect 450 70 485 75
rect 515 70 550 75
rect 390 60 435 70
rect 420 45 435 60
rect 395 40 435 45
rect 300 10 375 20
rect 390 30 435 40
rect 390 15 405 30
rect 420 15 435 30
rect 245 5 285 10
rect 305 5 370 10
rect 390 5 435 15
rect 250 0 285 5
rect 310 0 330 5
rect 345 0 365 5
rect 395 0 435 5
rect 450 65 490 70
rect 450 55 495 65
rect 450 0 465 55
rect 480 45 495 55
rect 510 60 555 70
rect 510 45 525 60
rect 540 45 555 60
rect 510 30 555 45
rect 510 15 525 30
rect 510 5 555 15
rect 515 0 555 5
<< end >>
