magic
tech sky130A
timestamp 1598774184
<< metal1 >>
rect 0 90 15 105
rect 0 75 20 90
rect 0 70 25 75
rect 5 65 25 70
rect 5 60 30 65
rect 10 55 30 60
rect 10 50 35 55
rect 15 45 35 50
rect 15 40 40 45
rect 20 35 40 40
rect 20 30 45 35
rect 25 15 45 30
rect 30 0 45 15
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
