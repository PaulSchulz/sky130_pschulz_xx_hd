magic
tech sky130A
timestamp 1598538767
<< metal1 >>
rect -725 675 -695 705
rect -725 645 -695 660
rect -710 585 -695 645
rect -725 575 -695 585
rect -725 570 -700 575
<< properties >>
string FIXED_BBOX 0 0 -130nm 1050nm
<< end >>
