magic
tech sky130A
timestamp 1598786878
<< metal1 >>
rect 0 0 30 30
<< properties >>
string FIXED_BBOX 0 -30 45 105
<< end >>
