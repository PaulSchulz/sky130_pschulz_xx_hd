magic
tech sky130A
timestamp 1598776905
<< metal1 >>
rect 0 70 30 75
rect 45 70 65 75
rect 0 65 70 70
rect 0 55 75 65
rect 0 0 15 55
rect 30 0 45 55
rect 60 0 75 55
<< properties >>
string FIXED_BBOX 0 -30 90 105
<< end >>
