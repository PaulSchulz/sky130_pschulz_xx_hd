magic
tech sky130A
timestamp 1598787399
<< metal1 >>
rect 0 45 30 75
rect 0 0 30 30
<< properties >>
string FIXED_BBOX 0 -30 45 105
<< end >>
