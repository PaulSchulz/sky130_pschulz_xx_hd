magic
tech sky130A
timestamp 1598786195
<< metal1 >>
rect 20 100 55 105
rect 15 95 60 100
rect 10 85 65 95
rect 10 80 25 85
rect 5 70 25 80
rect 50 70 65 85
rect 5 65 30 70
rect 10 60 35 65
rect 10 55 40 60
rect 10 50 45 55
rect 5 45 50 50
rect 0 40 55 45
rect 0 35 20 40
rect 35 35 60 40
rect 0 20 15 35
rect 40 30 65 35
rect 40 25 70 30
rect 40 20 75 25
rect 0 15 20 20
rect 35 15 75 20
rect 0 10 75 15
rect 5 5 75 10
rect 10 0 45 5
rect 60 0 75 5
<< properties >>
string FIXED_BBOX 0 -30 90 105
<< end >>
