magic
tech sky130A
timestamp 1598763351
<< metal1 >>
rect 10 100 45 105
rect 5 95 45 100
rect 0 85 45 95
rect 0 20 15 85
rect 0 10 45 20
rect 5 5 45 10
rect 10 0 45 5
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
