magic
tech sky130A
timestamp 1598777815
<< metal1 >>
rect 0 55 15 75
rect 30 55 45 75
rect 0 45 45 55
rect 5 30 40 45
rect 0 20 45 30
rect 0 0 15 20
rect 30 0 45 20
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
