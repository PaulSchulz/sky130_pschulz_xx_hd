magic
tech sky130A
timestamp 1598768855
<< metal1 >>
rect 10 100 45 105
rect 5 95 45 100
rect 0 85 45 95
rect 0 65 15 85
rect 0 60 35 65
rect 0 55 40 60
rect 5 50 45 55
rect 10 45 45 50
rect 30 20 45 45
rect 0 10 45 20
rect 0 5 40 10
rect 0 0 35 5
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
