magic
tech sky130A
timestamp 1598776260
<< metal1 >>
rect 0 75 30 105
rect 0 45 30 60
rect 15 15 30 45
rect 0 0 30 15
<< properties >>
string FIXED_BBOX 0 -30 45 105
<< end >>
