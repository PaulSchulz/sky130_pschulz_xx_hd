magic
tech sky130A
timestamp 1598777411
<< metal1 >>
rect 0 20 15 75
rect 30 20 45 75
rect 0 10 45 20
rect 5 5 45 10
rect 10 0 45 5
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
