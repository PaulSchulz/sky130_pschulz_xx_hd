magic
tech sky130A
timestamp 1598786008
<< metal1 >>
rect 15 75 30 105
rect 45 75 60 105
rect 0 60 75 75
rect 15 45 30 60
rect 45 45 60 60
rect 0 30 75 45
rect 15 0 30 30
rect 45 0 60 30
<< properties >>
string FIXED_BBOX 0 -30 90 105
<< end >>
