magic
tech sky130A
timestamp 1598786350
<< metal1 >>
rect 0 100 20 105
rect 0 95 25 100
rect 0 85 30 95
rect 15 20 30 85
rect 0 10 30 20
rect 0 5 25 10
rect 0 0 20 5
<< properties >>
string FIXED_BBOX 0 -30 45 105
<< end >>
