magic
tech sky130A
timestamp 1598786817
<< metal1 >>
rect 0 45 60 60
<< properties >>
string FIXED_BBOX 0 -30 75 105
<< end >>
