magic
tech sky130A
timestamp 1598775086
<< metal1 >>
rect 0 75 30 105
rect 0 60 15 75
<< properties >>
string FIXED_BBOX 0 -30 45 105
<< end >>
