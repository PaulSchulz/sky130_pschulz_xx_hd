magic
tech sky130A
timestamp 1598775974
<< metal1 >>
rect 20 100 45 105
rect 15 90 45 100
rect 15 75 30 90
rect 0 60 45 75
rect 15 0 30 60
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
