magic
tech sky130A
timestamp 1598784793
<< metal1 >>
rect 25 100 45 105
rect 20 95 45 100
rect 15 85 45 95
rect 15 70 30 85
rect 10 60 30 70
rect 0 45 25 60
rect 10 35 30 45
rect 15 20 30 35
rect 15 10 45 20
rect 20 5 45 10
rect 25 0 45 5
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
